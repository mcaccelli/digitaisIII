ataera.vhdl
